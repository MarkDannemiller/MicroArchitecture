
module coinCounter (
    
);
    
endmodule