//`include "debug_defs.v"

module top(
    input wire clk,                  // System clock signal that drives all pipeline stages
    input wire rst                   // Active-high reset signal to initialize all pipeline registers
);
    // ========================================================================
    // Pipeline Stage Signals and Registers - Detailed Description
    // ========================================================================
    /*
     * This RISC CPU implements a 4-stage pipeline:
     * 1. IF  (Instruction Fetch)    - Retrieves instruction from memory, calculates next PC
     * 2. DOF (Decode & Operand Fetch) - Decodes instruction, reads register file, prepares operands
     * 3. EX  (Execute)              - Performs ALU operations, memory access, branch calculation
     * 4. WB  (Write Back)           - Writes results back to register file
     * 
     * Each pipeline stage has its own dedicated module that performs specific operations.
     * Data flows between stages through pipeline registers that are updated on negative clock edges.
     * This prevents data hazards and ensures correct operation timing.
     */
    
    // Program Counter Registers - Track instruction execution across pipeline stages
    reg [31:0] PC;      // Current Program Counter for IF stage (points to current instruction)
    reg [31:0] PC_1;    // PC+1 value passed to DOF stage (for jump-and-link instructions)
    reg [31:0] PC_2;    // PC+2 value passed to EX and WB stages (for branch target calculation)
    
    // IF Stage output signals - Retrieved from Instruction Fetch module
    wire [31:0] IF_PC_next;     // Next PC value calculated by MuxC (based on branch/jump decisions)
    wire [31:0] IF_PC_plus_1;   // PC+1 from incrementer (sequential next instruction address)
    wire [31:0] IF_instruction; // Current instruction fetched from instruction memory
    
    // IF to DOF Pipeline Register - Passes fetched instruction to decode stage
    reg [31:0] IF_DOF_instruction; // Instruction register that holds fetched instruction for DOF stage
    
    // DOF Stage output signals - Generated by Decode & Operand Fetch module
    wire [31:0] DOF_A_data;         // Data read from register A (source register 1)
    wire [31:0] DOF_B_data;         // Data read from register B (source register 2)
    wire [31:0] DOF_BusA;           // Output from MuxA - selects between register A and PC+1
    wire [31:0] DOF_BusB;           // Output from MuxB - selects between register B and immediate value
    wire [31:0] DOF_extended_imm;   // Sign/zero-extended immediate value from instruction
    wire DOF_RW;                    // Register Write control signal - indicates if instruction writes to register
    wire DOF_MW;                    // Memory Write control signal - indicates if instruction writes to memory
    wire [1:0] DOF_MD;              // Memory Data select (2 bits) - selects source for register write data
    wire [1:0] DOF_BS;              // Branch Select control - determines branch type (no branch/conditional/register/direct)
    wire DOF_PS;                    // Program Select control - selects branch condition polarity (BZ vs BNZ)
    wire [4:0] DOF_FS;              // Function Select code - determines ALU operation
    wire [4:0] DOF_DR;              // Destination Register number - target register for write operations
    wire [4:0] DOF_SH;              // Shift amount field - for shift instructions (LSL, LSR)
    
    // DOF to EX Pipeline Registers - Pass decode output signals to execute stage
    reg [31:0] DOF_EX_BusA;           // Bus A value from DOF stage (first ALU operand)
    reg [31:0] DOF_EX_BusB;           // Bus B value from DOF stage (second ALU operand)
    reg [31:0] DOF_EX_extended_imm;   // Extended immediate value (for memory and branch address calculation)
    reg DOF_EX_RW;                    // Register Write control (pipelined to EX stage)
    reg [1:0] DOF_EX_MD;              // Memory Data select (pipelined to EX stage)
    reg DOF_EX_MW;                    // Memory Write control (pipelined to EX stage)
    reg [4:0] DOF_EX_FS;              // Function Select (pipelined to EX stage)
    reg [4:0] DOF_EX_DR;              // Destination Register (pipelined to EX stage)
    reg [4:0] DOF_EX_SH;              // Shift amount (pipelined to EX stage)
    reg [1:0] DOF_EX_BS;              // Branch Select (pipelined to EX stage)
    reg DOF_EX_PS;                    // Program Select (pipelined to EX stage)
    
    // EX Stage output signals - Generated by Execute module
    wire [31:0] EX_ALU_result;     // Result of ALU operation
    wire [31:0] EX_mem_data;       // Data read from memory (for load instructions)
    wire EX_Z;                     // Zero flag - set when ALU result is zero
    wire EX_V;                     // Overflow flag - set when arithmetic overflow occurs
    wire EX_N;                     // Negative flag - set when ALU result is negative (MSB=1)
    wire EX_C;                     // Carry flag - set when arithmetic carry/borrow occurs
    wire EX_N_xor_V;               // N XOR V condition - used for signed comparison (SLT)
    wire [31:0] EX_BrA;            // Calculated branch target address
    
    // EX to WB Pipeline Registers - Pass execute results to writeback stage
    reg [31:0] EX_WB_ALU_result;   // ALU result from EX stage (for register write operations)
    reg [31:0] EX_WB_mem_data;     // Memory data from EX stage (for load operations)
    reg EX_WB_N_xor_V;             // N XOR V condition (pipelined to WB stage for SLT)
    reg [1:0] EX_WB_MD;            // Memory Data select (pipelined to WB stage)
    reg EX_WB_RW;                  // Register Write control (pipelined to WB stage)
    reg [4:0] EX_WB_DR;            // Destination Register (pipelined to WB stage)
    
    // WB Stage output signals - Generated by Writeback module
    wire [31:0] WB_data;           // Final data to write to register file
    wire [4:0] WB_addr;            // Final register address to write to
    wire WB_en;                    // Final write enable signal for register file

    // ========================================================================
    // Pipeline Stage Module Instantiations
    // ========================================================================

    // IF Stage - Instruction Fetch
    /*
     * The IF stage fetches the next instruction from instruction memory
     * and calculates the next PC value based on branch/jump conditions.
     * 
     * Key operations:
     * - Fetches instruction at current PC from instruction memory
     * - Calculates PC+1 for sequential execution
     * - Selects next PC value based on branch/jump conditions
     */
    IF_stage if_stage(
        .clk(clk),                  // System clock
        .rst(rst),                  // Reset signal
        .PC(PC),                    // Current Program Counter (input to instruction memory)
        .BrA(EX_BrA),               // Branch target address (calculated in EX stage)
        .RAA(DOF_EX_BusA),          // Jump register address (for JMR - jump to register)
        .JMP(EX_BrA),               // Jump target address (for JMP - direct jump)
        .BS(DOF_EX_BS),             // Branch control from DOF (pipelined through EX)
        .PS(DOF_EX_PS),             // Program select from DOF (pipelined through EX)
        .Z(EX_Z),                   // Zero flag from EX stage (for conditional branches)
        .PC_next(IF_PC_next),       // Next PC value output (to update PC register)
        .PC_1(IF_PC_plus_1),        // PC+1 output (for sequential execution and JML)
        .instruction(IF_instruction) // Fetched instruction output
    );

    // DOF Stage - Decode & Operand Fetch
    /*
     * The DOF stage decodes the instruction, reads operands from the register file,
     * and generates control signals for subsequent pipeline stages.
     * 
     * Key operations:
     * - Decodes instruction opcode to generate control signals
     * - Reads source registers from register file
     * - Extends immediate values from instruction
     * - Selects operands for the ALU through MuxA and MuxB
     */
    DOF_stage dof_stage(
        .clk(clk),                   // System clock
        .rst(rst),                   // Reset signal
        .instruction(IF_DOF_instruction), // Instruction from IF stage (through pipeline register)
        .PC_1(PC_1),                 // PC+1 from pipeline register (for jump-and-link)
        .WB_data(WB_data),           // Write data from WB stage (for register write)
        .WB_addr(WB_addr),           // Write address from WB stage (register number)
        .WB_en(WB_en),               // Write enable from WB stage
        .A_data(DOF_A_data),         // Source register A data output
        .B_data(DOF_B_data),         // Source register B data output
        .BusA(DOF_BusA),             // MuxA output - first ALU operand
        .BusB(DOF_BusB),             // MuxB output - second ALU operand
        .extended_imm(DOF_extended_imm), // Extended immediate value
        .RW(DOF_RW),                 // Register Write control signal
        .MD(DOF_MD),                 // Memory Data select (2 bits for MuxD)
        .MW(DOF_MW),                 // Memory Write control signal
        .BS(DOF_BS),                 // Branch Select control signals
        .PS(DOF_PS),                 // Program Select (branch condition)
        .FS(DOF_FS),                 // Function Select (ALU operation)
        .DR(DOF_DR),                 // Destination Register number
        .SH(DOF_SH)                  // Shift amount field
    );

    // EX Stage - Execute
    /*
     * The EX stage performs the actual computation, memory access,
     * and branch target calculation.
     * 
     * Key operations:
     * - Performs ALU operations based on FS signal
     * - Accesses data memory for load/store operations
     * - Calculates branch target addresses
     * - Sets condition flags (Z, N, V, C) based on computation results
     */
    EX_stage ex_stage(
        .clk(clk),                   // System clock
        .rst(rst),                   // Reset signal
        .BusA(DOF_EX_BusA),          // First ALU operand from DOF stage
        .BusB(DOF_EX_BusB),          // Second ALU operand from DOF stage
        .extended_imm(DOF_EX_extended_imm), // Extended immediate for memory/branch address
        .PC_2(PC_2),                 // PC+2 from pipeline register (for branch calculation)
        .SH(DOF_EX_SH),              // Shift amount for barrel shifter operations
        .FS(DOF_EX_FS),              // Function Select code for ALU operation
        .MW(DOF_EX_MW),              // Memory Write control for store operations
        .ALU_result(EX_ALU_result),  // ALU computation result output
        .mem_data(EX_mem_data),      // Data read from memory (for load operations)
        .BrA(EX_BrA),                // Calculated branch target address output
        .N_xor_V(EX_N_xor_V),        // N XOR V condition for SLT instruction
        .Z(EX_Z),                    // Zero flag output
        .V(EX_V),                    // Overflow flag output
        .N(EX_N),                    // Negative flag output
        .C(EX_C)                     // Carry flag output
    );

    // WB Stage - Write Back
    /*
     * The WB stage selects and writes the computation result
     * back to the register file.
     * 
     * Key operations:
     * - Selects final write data from ALU result, memory data, or condition flag
     * - Generates final write enable signal based on RW control
     * - Passes final write address (destination register) to register file
     */
    WB_stage wb_stage(
        .ALU_result(EX_WB_ALU_result), // ALU result from EX stage
        .mem_data(EX_WB_mem_data),     // Memory data from EX stage
        .N_xor_V(EX_WB_N_xor_V),       // N XOR V condition for SLT instruction
        .MD(EX_WB_MD),                 // Memory Data select - chooses data source
        .RW(EX_WB_RW),                 // Register Write control from EX stage
        .DR(EX_WB_DR),                 // Destination Register from EX stage
        .WB_data(WB_data),             // Final data to write to register file
        .WB_addr(WB_addr),             // Final register address to write to
        .WB_en(WB_en)                  // Final write enable signal
    );

    // ========================================================================
    // Pipeline Registers Update Logic - Implements Pipelining Mechanism
    // ========================================================================
    
    // PC Pipeline Registers - Track instruction across pipeline stages
    /*
     * These registers track the PC values across pipeline stages.
     * They are updated on negative clock edge to ensure data is stable
     * when used by the next stage on positive clock edge.
     */
    always @(negedge clk or posedge rst) begin
        if (rst) begin
            // Initialize all PC registers to 0 on reset
            PC <= 32'h0;     // Starting address for program execution
            PC_1 <= 32'h0;   // Reset PC+1 register
            PC_2 <= 32'h0;   // Reset PC+2 register
        end
        else begin
            // Normal pipeline flow - PC values move through pipeline
            PC <= IF_PC_next;      // Update PC with next instruction address
            PC_1 <= IF_PC_plus_1;  // Update PC_1 with PC+1 value (for DOF stage)
            PC_2 <= PC_1;          // Update PC_2 with previous PC_1 (for EX stage)
        end
    end
    
    // IF to DOF Pipeline Register - Passes instruction to decode stage
    /*
     * This register passes the fetched instruction from IF to DOF stage.
     * Updated on negative edge to ensure instruction is stable for decoding.
     */
    always @(negedge clk or posedge rst) begin
        if (rst) begin
            // Reset instruction register to NOP
            IF_DOF_instruction <= 32'h0;
        end
        else begin
            // Latch the fetched instruction for decoding
            IF_DOF_instruction <= IF_instruction;
        end
    end
    
    // DOF to EX Pipeline Registers - Pass decode outputs to execute stage
    /*
     * These registers pass control signals and operands from DOF to EX stage.
     * They implement the pipeline structure that enables overlapped execution.
     */
    always @(negedge clk or posedge rst) begin
        if (rst) begin
            // Reset all pipeline registers to default values
            DOF_EX_BusA <= 32'h0;          // Reset operand A
            DOF_EX_BusB <= 32'h0;          // Reset operand B
            DOF_EX_extended_imm <= 32'h0;   // Reset extended immediate
            DOF_EX_RW <= 1'b0;             // Disable register write
            DOF_EX_MD <= 2'b00;            // Reset memory data select
            DOF_EX_MW <= 1'b0;             // Disable memory write
            DOF_EX_FS <= 5'h0;             // Reset function select (NOP)
            DOF_EX_DR <= 5'h0;             // Reset destination register (R0)
            DOF_EX_SH <= 5'h0;             // Reset shift amount
            DOF_EX_BS <= 2'b00;            // Reset branch select (no branch)
            DOF_EX_PS <= 1'b0;             // Reset program select
        end
        else begin
            // Pass DOF stage outputs to EX stage
            DOF_EX_BusA <= DOF_BusA;               // First ALU operand
            DOF_EX_BusB <= DOF_BusB;               // Second ALU operand
            DOF_EX_extended_imm <= DOF_extended_imm; // Extended immediate value
            DOF_EX_RW <= DOF_RW;                   // Register write control
            DOF_EX_MD <= DOF_MD;                   // Memory data select
            DOF_EX_MW <= DOF_MW;                   // Memory write control
            DOF_EX_FS <= DOF_FS;                   // Function select
            DOF_EX_DR <= DOF_DR;                   // Destination register
            DOF_EX_SH <= DOF_SH;                   // Shift amount
            DOF_EX_BS <= DOF_BS;                   // Branch select
            DOF_EX_PS <= DOF_PS;                   // Program select
        end
    end
    
    // EX to WB Pipeline Registers - Pass execute results to writeback stage
    /*
     * These registers pass computation results and control signals from EX to WB stage.
     * They enable pipelined execution where different instructions are at different stages.
     */
    always @(negedge clk or posedge rst) begin
        if (rst) begin
            // Reset all EX to WB pipeline registers
            EX_WB_ALU_result <= 32'h0;     // Reset ALU result
            EX_WB_mem_data <= 32'h0;       // Reset memory data
            EX_WB_N_xor_V <= 1'b0;         // Reset N XOR V condition
            EX_WB_RW <= 1'b0;              // Disable register write
            EX_WB_MD <= 2'b00;             // Reset memory data select
            EX_WB_DR <= 5'h0;              // Reset destination register
        end
        else begin
            // Pass EX stage outputs to WB stage
            EX_WB_ALU_result <= EX_ALU_result;  // ALU computation result
            EX_WB_mem_data <= EX_mem_data;      // Memory read data
            EX_WB_N_xor_V <= EX_N_xor_V;        // N XOR V condition for SLT
            EX_WB_RW <= DOF_EX_RW;              // Register write control
            EX_WB_MD <= DOF_EX_MD;              // Memory data select
            EX_WB_DR <= DOF_EX_DR;              // Destination register
            
            // Enhanced debug output for tracking register write through pipeline
            if (`DEBUG_PIPE) begin
                $display("PIPELINE DEBUG: DOF_RW=%b, DOF_EX_RW=%b -> EX_WB_RW=%b", 
                         DOF_RW, DOF_EX_RW, EX_WB_RW);
                $display("PIPELINE DEBUG: DR Path: DOF_DR=%d -> DOF_EX_DR=%d -> EX_WB_DR=%d", 
                         DOF_DR, DOF_EX_DR, DOF_EX_DR);
                $display("PIPELINE DEBUG: ALU_result=%h for instruction at PC=%h", 
                         EX_ALU_result, PC_2);
                $display("PIPELINE DEBUG: WB_data=%h, WB_addr=%d, WB_en=%b", 
                         WB_data, WB_addr, WB_en);
            end
        end
    end

    // Add debug output for instruction execution
    always @(posedge clk) begin
        if (!rst && `DEBUG_PIPE) begin
            $display("INSTRUCTION DEBUG: PC=%h, Instruction=%h", PC, IF_instruction);
            $display("INSTRUCTION DEBUG: Opcode=%b, DR=%d, SA=%d, SB=%d", 
                     IF_instruction[31:25], IF_instruction[24:20], 
                     IF_instruction[19:15], IF_instruction[14:10]);
        end
    end

    // Add debug output for register file updates
    always @(posedge clk) begin
        if (!rst && `DEBUG_PIPE && WB_en) begin
            $display("REGISTER DEBUG: Writing %h to R%d", WB_data, WB_addr);
        end
    end

endmodule
